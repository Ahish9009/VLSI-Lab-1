
module norGate(x, op);
input x;
output op;
assign op = ~(x);
endmodule
