
module notGate(x, op);
input x;
output op;
assign op = ~(x);
endmodule
